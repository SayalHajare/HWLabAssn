// Design a 16*4 mux from using 4*2 mux.
// Input consists of two arrays:
//          a. Data consisting of an array of size 16.
//          b. Select lines consisting of an array of size 4.
// Implement 4*2 mux in Verilog and then call its module within the module for 16*4 mux.
// Write test bench to simulate the behavior of the code.